module MinerBitMap (
    input   logic        clk,
    input   logic        resetN,
    input   logic [10:0] offsetX,
    input   logic [10:0] offsetY,
    input   logic        InsideRectangle,

    output logic        drawingRequest,
    output logic [7:0]  RGBout
);

    localparam logic [7:0] TRANSPARENT_ENCODING = 8'h72; 
    
    localparam int OBJECT_WIDTH_X = 128;
    localparam int OBJECT_HEIGHT_Y = 128;
	 
	 
    logic [0:OBJECT_HEIGHT_Y-1][0:OBJECT_WIDTH_X-1][7:0] object_colors = {
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h71,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'hF5,8'hF8,8'hF8,8'hF8,8'hF8,8'hF9,8'h20,8'h00,8'h00,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFD,8'h84,8'hF8,8'hF8,8'h00,8'h20,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h64,8'hFD,8'hFD,8'hFD,8'hFD,8'hFD,8'hF8,8'hF8,8'hFD,8'h20,8'hFC,8'hFD,8'hF5,8'h00,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h92,8'h00,8'hF8,8'hFD,8'hFD,8'hFD,8'hFD,8'hF8,8'hFC,8'hFD,8'h20,8'hF4,8'hFC,8'hFD,8'hFD,8'hFD,8'h20,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'hF9,8'hF8,8'hFD,8'hFF,8'hFF,8'hFF,8'hF8,8'hFC,8'hFC,8'h00,8'h60,8'hFC,8'hFD,8'hFD,8'hFD,8'hFC,8'hB1,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'hF8,8'hF4,8'hF8,8'hFC,8'hFF,8'hF8,8'hF8,8'hFC,8'hFC,8'hD0,8'h60,8'hF8,8'hFC,8'hFC,8'hFC,8'hFC,8'hF9,8'hF9,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'hD0,8'hF4,8'hF4,8'hF8,8'hF8,8'hFE,8'hF8,8'hF8,8'hF8,8'hF8,8'hAC,8'h60,8'hF8,8'hF8,8'hF8,8'hF8,8'hFC,8'hF8,8'hF4,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'hD0,8'hF4,8'hF4,8'hF4,8'hF4,8'hF8,8'hF4,8'hF4,8'hF4,8'hF4,8'hAC,8'h84,8'h20,8'h20,8'h20,8'hF0,8'hFC,8'hF8,8'hF4,8'h00,8'h04,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h00,8'h8C,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'h84,8'h64,8'hF8,8'hFC,8'h8C,8'hD0,8'hF4,8'hF8,8'hF0,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h92,8'h64,8'h64,8'h84,8'hD0,8'hD0,8'hD0,8'hD0,8'hF0,8'hD0,8'hF0,8'hF0,8'hF0,8'hD0,8'hD0,8'hD0,8'h20,8'hF4,8'hF4,8'h84,8'hF4,8'h84,8'hF5,8'hF0,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h04,8'h00,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF5,8'hF5,8'hF5,8'hF5,8'hF5,8'h64,8'hF8,8'hF9,8'h00,8'hB1,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'hB1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'hF9,8'h84,8'hF9,8'hAC,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'h00,8'hF5,8'hD1,8'hD5,8'hD6,8'hF1,8'hF1,8'hF1,8'hF1,8'h20,8'h20,8'h20,8'hD5,8'hF1,8'hF1,8'hB1,8'h00,8'h00,8'h00,8'h00,8'hF4,8'hF5,8'hAC,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h92,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFA,8'hFA,8'hFA,8'hFA,8'h00,8'h00,8'h00,8'h00,8'hFA,8'hF9,8'hD1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'hD1,8'h00,8'h71,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hFA,8'hFA,8'hFA,8'hFE,8'hFA,8'hFF,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hB1,8'h20,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hF6,8'hFF,8'h00,8'h24,8'hFF,8'hFE,8'hFF,8'hFF,8'hFF,8'h00,8'hFF,8'h20,8'hFF,8'hFF,8'h91,8'h20,8'h20,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h00,8'hF6,8'hFF,8'h00,8'h24,8'hFF,8'hFE,8'hFF,8'hFF,8'hFF,8'h00,8'h6D,8'h20,8'hFF,8'hFF,8'h91,8'h20,8'h91,8'hFF,8'hFE,8'hFE,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h92,8'h00,8'hF6,8'hFF,8'h00,8'h00,8'h00,8'hFE,8'hFE,8'hFF,8'hFF,8'h00,8'h00,8'h24,8'hFF,8'hFF,8'h91,8'h20,8'hFF,8'h00,8'h20,8'hF9,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h00,8'hF6,8'hF6,8'hFF,8'hFF,8'h00,8'hFE,8'hFE,8'hFE,8'hB1,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'h20,8'h20,8'h64,8'h20,8'h60,8'hD5,8'hF9,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'hF5,8'hFE,8'h00,8'h20,8'h00,8'hD1,8'hD5,8'hD1,8'h00,8'h20,8'h20,8'h20,8'hFF,8'hFF,8'h20,8'h20,8'hFA,8'h20,8'h84,8'hFE,8'hFE,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'hF6,8'h20,8'h20,8'h20,8'h20,8'h00,8'h00,8'h00,8'h20,8'h20,8'h20,8'h20,8'h00,8'hFF,8'h20,8'h20,8'h20,8'h20,8'hFE,8'hFA,8'h00,8'h24,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'h20,8'h20,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h20,8'h20,8'h00,8'h20,8'h20,8'h20,8'h00,8'h00,8'h00,8'h25,8'h2D,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h20,8'h20,8'h20,8'h00,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h20,8'h20,8'h20,8'h20,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h20,8'h20,8'h20,8'h20,8'h60,8'h60,8'h60,8'h60,8'h64,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h00,8'h71,8'h72,8'h71,8'h71,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h92,8'h00,8'h20,8'h20,8'h20,8'h20,8'h60,8'h84,8'h84,8'h84,8'h84,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h00,8'h71,8'h92,8'h00,8'h00,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h92,8'h92,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h00,8'h00,8'hD1,8'h00,8'h00,8'h76,8'h77,8'h96,8'h00,8'h00,8'h00,8'h00,8'h24,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h6D,8'h00,8'h00,8'h00,8'h00,8'h76,8'h76,8'h00,8'h00,8'h00,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h00,8'h00,8'h20,8'hD1,8'hD1,8'h00,8'h77,8'h76,8'h04,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFA,8'h00,8'h00,8'h00,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'hFE,8'hB1,8'h00,8'h76,8'h76,8'h00,8'h20,8'h20,8'h00,8'h00,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h00,8'h85,8'h8D,8'hB1,8'hD5,8'h72,8'h76,8'h76,8'h00,8'hF0,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hFE,8'hFE,8'hFE,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h92,8'h00,8'hF9,8'hFE,8'hF4,8'h84,8'h2D,8'h76,8'h76,8'h00,8'hC4,8'hEC,8'h20,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'hF1,8'hF5,8'hD1,8'h00,8'h76,8'h76,8'h76,8'h20,8'hF4,8'hF4,8'hF4,8'hF4,8'hFE,8'hF4,8'hF4,8'hF4,8'hF9,8'hFE,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h00,8'hFA,8'hF4,8'hF4,8'hF4,8'h64,8'h2D,8'h76,8'h76,8'h00,8'hEC,8'hEC,8'hC4,8'hA4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hF1,8'hF1,8'hF5,8'h60,8'h20,8'h00,8'h72,8'h76,8'h76,8'h20,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hFE,8'h20,8'h00,8'h2D,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'hFE,8'hF4,8'hF4,8'hF4,8'hF4,8'h64,8'h2D,8'h76,8'h76,8'h00,8'hEC,8'hEC,8'h00,8'h00,8'hD1,8'hF1,8'hF1,8'hF1,8'hF1,8'hF1,8'hF1,8'hD1,8'h00,8'h00,8'hF0,8'hF5,8'h00,8'h72,8'h32,8'h72,8'h20,8'hF0,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF9,8'hFE,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h2D,8'h00,8'hFD,8'hF4,8'hF4,8'hF4,8'hF4,8'h64,8'h2D,8'h76,8'h76,8'h00,8'hF0,8'hF0,8'hC4,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h00,8'hF0,8'hF4,8'hF5,8'h00,8'h72,8'h32,8'h32,8'h20,8'hF0,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF9,8'hFE,8'h00,8'h71,8'h2D,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hFE,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'h64,8'h2D,8'h76,8'h76,8'h00,8'hF0,8'hF0,8'hC4,8'hA4,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'hF4,8'hF0,8'hF4,8'h00,8'h32,8'h32,8'h32,8'h20,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF9,8'h00,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'hFD,8'hF4,8'hF4,8'hF4,8'hF4,8'hF0,8'h64,8'h2D,8'h76,8'h76,8'h00,8'hF0,8'hF0,8'hF0,8'hEC,8'hEC,8'hEC,8'hCC,8'hCC,8'hC4,8'hCC,8'hF0,8'hF0,8'hF4,8'hF4,8'hF4,8'hCC,8'h00,8'h2D,8'h2E,8'h2D,8'h20,8'hF4,8'hF4,8'hF0,8'hF0,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hFD,8'h00,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h00,8'h00,8'hFD,8'hF4,8'hF4,8'hF4,8'hC4,8'hA4,8'h84,8'h25,8'h2D,8'h2D,8'h00,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF4,8'hF4,8'hF0,8'hF0,8'hEC,8'h00,8'h2D,8'h2D,8'h2D,8'h20,8'hEC,8'hC4,8'hEC,8'hF0,8'hF0,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF5,8'h64,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h00,8'hFD,8'hF4,8'hF4,8'hF4,8'hF4,8'hC4,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'hEC,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF4,8'hEC,8'h60,8'h00,8'h00,8'h00,8'h00,8'h20,8'hEC,8'hC4,8'hF0,8'hF0,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'h84,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h71,8'h25,8'h00,8'hFD,8'hF4,8'hF4,8'hF4,8'hF4,8'hCC,8'h20,8'hD5,8'hF5,8'hF5,8'hF5,8'h00,8'h20,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h20,8'h00,8'hF5,8'hF9,8'hF9,8'hF9,8'h20,8'hCC,8'hA4,8'hC4,8'hF0,8'hF4,8'hF4,8'hF0,8'hF4,8'hF4,8'hF4,8'hF4,8'hF4,8'h20,8'hD5,8'hFE,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h00,8'hFE,8'hF5,8'hF0,8'hF4,8'hF0,8'hF4,8'hCC,8'h20,8'hAC,8'h84,8'h84,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hF4,8'h84,8'h84,8'hF4,8'h20,8'hCC,8'h84,8'hEC,8'hC4,8'hF0,8'hF4,8'h80,8'hF0,8'hF0,8'hF5,8'h20,8'hFE,8'hFE,8'hFE,8'hFD,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h20,8'hF9,8'hF9,8'h60,8'hF0,8'hF4,8'hF0,8'hCC,8'h20,8'hAC,8'h60,8'h84,8'hF0,8'h00,8'h2D,8'h2D,8'h72,8'h72,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h00,8'hF4,8'h60,8'h84,8'hF4,8'h20,8'hC4,8'h84,8'hEC,8'hEC,8'hC4,8'hF0,8'hF0,8'hF1,8'h20,8'hFE,8'hFE,8'hFD,8'hFD,8'hF9,8'hF9,8'h20,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h6D,8'h20,8'hF5,8'hF9,8'hF9,8'hFE,8'h60,8'hF0,8'hC4,8'h20,8'h8D,8'hAC,8'hAC,8'hB0,8'h00,8'h2D,8'h2D,8'h72,8'h72,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h00,8'h8C,8'hAC,8'hAC,8'hAC,8'h20,8'hCC,8'h00,8'hC4,8'hEC,8'hEC,8'hA4,8'h20,8'hF9,8'hFE,8'hFE,8'hF9,8'hF9,8'hF9,8'hF5,8'h20,8'h20,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h00,8'hF5,8'hF5,8'hF9,8'hF9,8'hF0,8'h20,8'h84,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'hC4,8'h00,8'hC4,8'h20,8'h84,8'hF5,8'hF5,8'hF9,8'hF9,8'hF9,8'hF5,8'hF9,8'h20,8'h20,8'hFA,8'h00,8'h00,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h00,8'h8D,8'h20,8'hF9,8'hF5,8'hF0,8'hF0,8'hCD,8'h20,8'h00,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2E,8'h25,8'h25,8'h00,8'hC4,8'hC4,8'hC4,8'h00,8'h84,8'hCC,8'hF1,8'hF5,8'hF1,8'hF5,8'hF5,8'hB1,8'h20,8'hB1,8'hFE,8'hFF,8'hFF,8'h00,8'h00,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'hFE,8'hD1,8'h20,8'hD1,8'hF0,8'hF0,8'hCC,8'hF0,8'h00,8'h05,8'h2D,8'h2D,8'h2D,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h76,8'h76,8'h76,8'h32,8'h72,8'h72,8'h00,8'hF0,8'hF0,8'hCC,8'h00,8'hCC,8'hCC,8'hCC,8'hF1,8'hF1,8'h20,8'h00,8'hF5,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h92,8'h00,8'hFE,8'hFE,8'hF5,8'hD5,8'h00,8'hF1,8'hEC,8'hAC,8'h00,8'h04,8'h2D,8'h2D,8'h2D,8'h00,8'h76,8'h76,8'h9B,8'h9F,8'h9F,8'hBF,8'hBF,8'hBF,8'hBF,8'hBF,8'hFF,8'h00,8'h76,8'h76,8'h76,8'h72,8'h72,8'h00,8'hF0,8'hF0,8'hF0,8'hA4,8'h20,8'hAD,8'hCD,8'h20,8'h20,8'hFA,8'hFE,8'hFE,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hDA,8'hDA,8'hFE,8'hFE,8'hFE,8'hFE,8'hD1,8'hD1,8'h20,8'h60,8'h00,8'h05,8'h2D,8'h2D,8'h2D,8'h00,8'h36,8'h76,8'h7B,8'h7F,8'h7F,8'h7F,8'h7F,8'h7F,8'h7F,8'h7F,8'hFF,8'h00,8'h76,8'h76,8'h76,8'h76,8'h72,8'h00,8'hF0,8'hF0,8'hF0,8'hC4,8'h20,8'h20,8'h20,8'hCD,8'hCD,8'hF5,8'hF5,8'hF5,8'hF5,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h00,8'hFF,8'hFF,8'hFF,8'hF5,8'hF5,8'hFE,8'hFF,8'hD1,8'hD1,8'hB1,8'h00,8'h05,8'h2D,8'h2D,8'h2D,8'h00,8'h36,8'h76,8'h7B,8'h7B,8'h7F,8'h7F,8'h7F,8'h7F,8'h7F,8'h7F,8'hFF,8'h00,8'h76,8'h76,8'h76,8'h76,8'h72,8'h00,8'h00,8'h84,8'hF9,8'hCC,8'hA4,8'h20,8'h60,8'h84,8'h8C,8'hF5,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hFF,8'hFF,8'hFE,8'hFF,8'hFA,8'hF1,8'hD1,8'hD1,8'hCD,8'hCD,8'h00,8'h05,8'h2D,8'h2D,8'h2D,8'h00,8'h36,8'h76,8'h7B,8'h7B,8'h7B,8'h7F,8'h7B,8'h7F,8'h7F,8'h7F,8'hFF,8'h00,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h00,8'h60,8'hEC,8'hCC,8'hC4,8'h20,8'h00,8'hF5,8'hF5,8'hFE,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h25,8'h00,8'hFF,8'hFE,8'hFE,8'hFE,8'hFF,8'hFF,8'hFA,8'hF1,8'hD1,8'hCD,8'h00,8'h04,8'h2D,8'h2D,8'h2D,8'h00,8'h76,8'h76,8'h7B,8'h7F,8'h7F,8'h7F,8'h7F,8'h7F,8'h7F,8'h7F,8'hFF,8'h00,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h00,8'h80,8'hEC,8'hE4,8'hCC,8'h20,8'h00,8'hF5,8'hF5,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF5,8'hF5,8'hF5,8'hF5,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hFF,8'hFF,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF9,8'hF5,8'hD1,8'hCD,8'h00,8'h04,8'h2D,8'h2D,8'h2D,8'h00,8'h76,8'h76,8'hBF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h00,8'h80,8'hC4,8'hCC,8'h20,8'h00,8'h00,8'hF5,8'hF5,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF5,8'hF5,8'hF6,8'hF5,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'hFF,8'hFF,8'hFE,8'hFE,8'hFE,8'hFF,8'hFE,8'hF5,8'hF5,8'hD1,8'hCD,8'h00,8'h04,8'h2D,8'h2D,8'h2D,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h00,8'h64,8'hAC,8'hCC,8'h20,8'h00,8'h00,8'hF5,8'hF5,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,8'hF5,8'hF5,8'h8C,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h00,8'hFF,8'hFF,8'hFF,8'hFE,8'hFE,8'hFE,8'hFE,8'hF6,8'hF5,8'hCD,8'hCD,8'h00,8'h04,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h72,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h00,8'h00,8'hC4,8'h20,8'h00,8'h00,8'hF5,8'hF5,8'hFE,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,8'hFF,8'hFE,8'hFA,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h00,8'hFF,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'hF6,8'hD1,8'h00,8'h00,8'h05,8'h2D,8'h2D,8'h2D,8'h32,8'h2E,8'h72,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h2D,8'h00,8'h00,8'h00,8'h00,8'hF5,8'hF5,8'hFE,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,8'hFE,8'hFE,8'hFE,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hFE,8'hFE,8'hFE,8'hFF,8'hFF,8'hFE,8'hFE,8'hF5,8'hF6,8'hD1,8'h00,8'h00,8'h00,8'h05,8'h05,8'h05,8'h05,8'h05,8'h2D,8'h2D,8'h2E,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2E,8'h2E,8'h32,8'hBF,8'h9F,8'h9F,8'h2D,8'h2D,8'h32,8'h32,8'h25,8'h25,8'h2D,8'h00,8'h00,8'h00,8'hF5,8'hF5,8'hFE,8'hFF,8'hFF,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFF,8'hFF,8'hFE,8'hF5,8'hF5,8'h00,8'h00,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h2E,8'h2E,8'h76,8'h76,8'h76,8'h01,8'h76,8'h05,8'h76,8'h76,8'h76,8'h76,8'h76,8'h96,8'hBF,8'hBF,8'h2D,8'h76,8'h76,8'h76,8'h2E,8'h2D,8'h2D,8'h00,8'h00,8'h00,8'hF5,8'hF5,8'hFE,8'hFF,8'hFF,8'hFF,8'hFE,8'hFE,8'hFE,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'hF5,8'hF6,8'hF5,8'h00,8'h72,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h01,8'h76,8'h05,8'h76,8'h76,8'h76,8'h76,8'h76,8'h25,8'h25,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h2E,8'h2D,8'h2D,8'h00,8'h00,8'h00,8'hF5,8'hF5,8'hFE,8'hFF,8'hFE,8'hFF,8'hFE,8'hFE,8'hFE,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'hF5,8'h00,8'h00,8'h00,8'h71,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h05,8'h05,8'h2D,8'h2D,8'h2D,8'h00,8'h76,8'h05,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2E,8'h2E,8'h2D,8'h2D,8'h00,8'h00,8'h00,8'h00,8'hF5,8'hF5,8'hFF,8'hFF,8'hFE,8'hFE,8'hFA,8'hF6,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'hF5,8'hF6,8'h00,8'h25,8'h71,8'h72,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h2E,8'h72,8'h76,8'h76,8'h05,8'h76,8'h05,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2E,8'h2D,8'h00,8'hFA,8'h00,8'h00,8'hF5,8'hF5,8'hFE,8'hFE,8'hFE,8'hFE,8'hFA,8'hF6,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'h20,8'h00,8'h00,8'h72,8'h72,8'h72,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h2E,8'h2D,8'h76,8'h76,8'h76,8'h05,8'h76,8'h05,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h00,8'h00,8'h00,8'hF1,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h04,8'h00,8'hFF,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h05,8'h76,8'h05,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h00,8'h00,8'h00,8'hF1,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFF,8'hFE,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'h20,8'h00,8'h72,8'h72,8'h00,8'h25,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h05,8'h76,8'h05,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h00,8'h00,8'h00,8'hD1,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'hFE,8'hFE,8'hF5,8'h20,8'h00,8'h71,8'h71,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h01,8'h2D,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h00,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'hF5,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'h00,8'hFE,8'hFE,8'hFE,8'hD5,8'hAD,8'hFE,8'hFE,8'hF5,8'h20,8'h00,8'h00,8'h00,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h00,8'h2D,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h00,8'h00,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hFE,8'hF5,8'hF5,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h20,8'hFE,8'hFE,8'hFE,8'hF5,8'h00,8'hB1,8'hF6,8'hF5,8'h00,8'h00,8'h00,8'h00,8'h2D,8'h72,8'h76,8'h76,8'h76,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h00,8'h2D,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h00,8'h00,8'hF5,8'hF5,8'hF5,8'hF6,8'hFE,8'hFE,8'hFE,8'hFA,8'hF5,8'hF5,8'h24,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h04,8'h00,8'hF5,8'hFE,8'hFE,8'hFE,8'hF5,8'h00,8'hF6,8'hF5,8'h00,8'h00,8'h00,8'h00,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h72,8'h72,8'h2D,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h00,8'h00,8'h20,8'hF1,8'hF5,8'hF5,8'hF5,8'hF5,8'hF5,8'hF5,8'h20,8'h00,8'h24,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h71,8'h00,8'hF5,8'hFE,8'hFE,8'hF5,8'hF1,8'h20,8'h00,8'h00,8'h72,8'h00,8'h2D,8'h72,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h72,8'h2D,8'h2D,8'h6D,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2D,8'h2D,8'h2D,8'h00,8'hD1,8'hD1,8'hD1,8'hD1,8'hD1,8'h20,8'h20,8'h00,8'h00,8'h04,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'hAD,8'hF5,8'hF1,8'hF1,8'h20,8'h00,8'h00,8'h71,8'h00,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h72,8'h2D,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h72,8'h2D,8'h00,8'h00,8'h60,8'hD1,8'hD1,8'hD1,8'h20,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h25,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h71,8'h72,8'h71,8'h00,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h72,8'h2D,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2D,8'h76,8'h76,8'h76,8'h76,8'h76,8'h9B,8'h9B,8'h9B,8'h9B,8'h2D,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h71,8'h72,8'h72,8'h92,8'h72,8'h72,8'h71,8'h00,8'h2D,8'h32,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h72,8'h2D,8'h25,8'h25,8'h00,8'h00,8'h6D,8'h6D,8'h71,8'h00,8'h00,8'h2D,8'h72,8'h76,8'h76,8'h77,8'h9F,8'h9F,8'h9F,8'h9B,8'h2D,8'h2D,8'h00,8'h24,8'h6D,8'h6D,8'h6D,8'h6D,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h71,8'h72,8'h72,8'h71,8'h00,8'h76,8'h7B,8'h9B,8'h76,8'h76,8'h76,8'h76,8'h76,8'h72,8'h2D,8'h25,8'h25,8'h00,8'h00,8'h72,8'h72,8'h72,8'h00,8'h00,8'h25,8'h72,8'h72,8'h76,8'h76,8'h7B,8'h9F,8'h7B,8'h9B,8'h76,8'h2D,8'h00,8'h04,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h71,8'h71,8'h00,8'h76,8'h7B,8'h9B,8'h76,8'h76,8'h76,8'h2D,8'h2D,8'h2D,8'h2D,8'h00,8'h00,8'h00,8'h6D,8'h71,8'h72,8'h72,8'h72,8'h00,8'h25,8'h72,8'h72,8'h76,8'h76,8'h7B,8'h7B,8'h7B,8'h9B,8'h9B,8'h76,8'h00,8'h04,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h00,8'h72,8'h32,8'h2D,8'h2D,8'h76,8'h76,8'h76,8'h2D,8'h2D,8'h2D,8'h2D,8'h00,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h00,8'h25,8'h72,8'h72,8'h72,8'h76,8'h7B,8'h7B,8'h7B,8'h7B,8'h9B,8'h76,8'h00,8'h04,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h6D,8'h2D,8'h2D,8'h2D,8'h32,8'h32,8'h32,8'h2D,8'h2D,8'h2D,8'h2D,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h25,8'h2D,8'h2D,8'h32,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h72,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h2E,8'h32,8'h2E,8'h72,8'h72,8'h2D,8'h25,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'h00,8'h25,8'h25,8'h2D,8'h72,8'h32,8'h72,8'h72,8'h72,8'h72,8'h76,8'h76,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h25,8'h2D,8'h2D,8'h72,8'h72,8'h2D,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h72,8'h2D,8'h2D,8'h2D,8'h72,8'h76,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h25,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h72,8'h72,8'h2D,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h72,8'h2D,8'h2D,8'h2D,8'h72,8'h76,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'h00,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h25,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2E,8'h72,8'h2D,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h72,8'h76,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hF9,8'hFD,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h25,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2E,8'h72,8'h2D,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h72,8'h72,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h04,8'hCC,8'hF0,8'hFC,8'hF8,8'h00,8'h71,8'h71,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h2D,8'h25,8'h2D,8'h2D,8'h2D,8'h2D,8'h2D,8'h25,8'h25,8'h25,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h2D,8'h2D,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h25,8'hCC,8'hCC,8'hF8,8'hF4,8'h00,8'h00,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h25,8'h2D,8'h25,8'h2D,8'h2D,8'h25,8'h25,8'h25,8'h25,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h2D,8'h2D,8'h00,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h04,8'h24,8'hAC,8'hAC,8'h84,8'h60,8'hF0,8'hF0,8'hFD,8'hF9,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h00,8'h6D,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h25,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h2D,8'h2D,8'h00,8'h00,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h20,8'hB0,8'h64,8'h84,8'h20,8'hF9,8'h20,8'hF0,8'hF0,8'hF4,8'hF4,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h00,8'h84,8'h8D,8'h8D,8'h8D,8'h84,8'h84,8'h84,8'h84,8'h84,8'h65,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h85,8'h85,8'h85,8'h8D,8'h8D,8'hAD,8'hB1,8'hB1,8'hB1,8'hB1,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'hAC,8'hF0,8'hA4,8'hF0,8'hB0,8'hB1,8'hF8,8'hF8,8'h20,8'h84,8'hF4,8'hF0,8'h20,8'h00,8'h6D,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h00,8'h00,8'h64,8'h64,8'h64,8'h64,8'h84,8'h64,8'h60,8'h60,8'h60,8'h60,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h64,8'h60,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8C,8'h8C,8'hAD,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'hAC,8'hAC,8'h84,8'hF0,8'hF0,8'hD0,8'hF0,8'hF4,8'hF4,8'h20,8'hF4,8'hF4,8'h20,8'h20,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h25,8'h00,8'h00,8'h00,8'h00,8'h20,8'h20,8'h20,8'h20,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h20,8'h20,8'h20,8'h00,8'h00,8'h64,8'h64,8'h00,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'hAC,8'hA4,8'hA4,8'hCC,8'hD0,8'h84,8'hCC,8'hCC,8'hF0,8'h84,8'hAC,8'hAC,8'h00,8'hF9,8'hF8,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h2D,8'h00,8'h20,8'h20,8'h20,8'h20,8'h60,8'h60,8'h60,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h20,8'h60,8'h20,8'h20,8'h00,8'h00,8'h20,8'h00,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h64,8'hA4,8'h84,8'hAC,8'hAC,8'h84,8'hCC,8'hCC,8'hA4,8'h64,8'h00,8'h84,8'h20,8'hEC,8'hF0,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h00,8'h00,8'h64,8'h20,8'h00,8'h20,8'h60,8'h60,8'h60,8'h00,8'h71,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'h20,8'h60,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8D,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h6D,8'hAC,8'hF0,8'hCC,8'h20,8'h64,8'hA4,8'h8C,8'h64,8'hA4,8'hA4,8'h64,8'hAC,8'hF8,8'h20,8'h20,8'hEC,8'hF0,8'h00,8'h71,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h84,8'h8C,8'h20,8'h64,8'h20,8'h60,8'h60,8'h60,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'h20,8'h60,8'h20,8'h20,8'h00,8'h00,8'h00,8'h00,8'h20,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h92,8'h92,8'h00,8'hCC,8'hCC,8'hA4,8'hA4,8'h00,8'h20,8'hF4,8'h20,8'h84,8'h64,8'hAC,8'hF0,8'hF0,8'hF0,8'h00,8'hCC,8'h84,8'hD1,8'h20,8'h04,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h20,8'hCC,8'hCC,8'hCC,8'hCC,8'hAC,8'hAC,8'h60,8'h20,8'h84,8'h84,8'h60,8'h20,8'h60,8'h60,8'h60,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h00,8'h20,8'h60,8'h00,8'h84,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hF0,8'hD0,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h60,8'h20,8'h20,8'h20,8'h20,8'hF0,8'hF4,8'hF0,8'h00,8'h20,8'hAC,8'hF0,8'hCC,8'hA4,8'h00,8'h00,8'hD0,8'hCC,8'hF5,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h84,8'hF1,8'hF1,8'hF1,8'hF5,8'hCC,8'hCC,8'h84,8'h64,8'h64,8'h60,8'h60,8'h60,8'h20,8'h00,8'h00,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'h20,8'h20,8'h20,8'h84,8'hA4,8'hA4,8'hA4,8'hA4,8'hA4,8'hA4,8'hCC,8'h00,8'h92,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'hCC,8'hF4,8'h60,8'hF0,8'hD0,8'hA4,8'h20,8'hA4,8'hCC,8'hCC,8'hAC,8'h8C,8'h84,8'hA4,8'hA4,8'h84,8'h84,8'h20,8'hF0,8'hAC,8'hCC,8'hF4,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h25,8'h00,8'h00,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'h00,8'h20,8'h20,8'h84,8'h84,8'hA4,8'hA4,8'hA4,8'hA4,8'hA4,8'hCC,8'h20,8'h00,8'h00,8'h72,8'h72,8'h72,8'h00,8'hA4,8'hAC,8'hAC,8'h60,8'hD0,8'hAC,8'h20,8'hF5,8'h20,8'hA4,8'hA4,8'h84,8'h84,8'h20,8'h84,8'h20,8'h20,8'h20,8'h20,8'hA4,8'hAC,8'h84,8'h60,8'h64,8'h00,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h2D,8'h00,8'h00,8'h20,8'h20,8'h20,8'h60,8'h60,8'h60,8'h60,8'h60,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h00,8'h00,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h00,8'h00,8'h00,8'h20,8'h60,8'h60,8'h64,8'h64,8'h64,8'h64,8'h84,8'h84,8'h84,8'h00,8'h00,8'h72,8'h72,8'h72,8'h00,8'hA4,8'hA4,8'h00,8'hAC,8'hA4,8'hAC,8'hAC,8'hF4,8'hF0,8'h20,8'h20,8'h20,8'hD0,8'hF4,8'h20,8'h00,8'hCC,8'h20,8'h00,8'h84,8'h20,8'h84,8'hEC,8'hCC,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h6D,8'h00,8'h00,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h64,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h00,8'h00,8'h71,8'h72,8'h71,8'h00,8'h84,8'h20,8'h84,8'h84,8'h84,8'h8C,8'h8C,8'h84,8'hCC,8'hA4,8'h00,8'h84,8'hA4,8'hAC,8'hCC,8'h00,8'hA4,8'hA4,8'h20,8'h64,8'h60,8'h84,8'hA4,8'hA4,8'h00,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h92,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h71,8'h71,8'h71,8'h71,8'h72,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h71,8'h72,8'h71,8'h71,8'h71,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h71,8'h71,8'h72,8'h72,8'h71,8'h71,8'h72,8'h71,8'h71,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h71,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'hDB,8'hDB,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'hDB,8'hDB,8'hDB,8'hDB,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'hDB,8'hDB,8'hDA,8'hDA,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'hDB,8'hDB,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h71,8'h72,8'h72,8'h72,8'h71,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h71,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h71,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72}
};



always_ff @(posedge clk or negedge resetN) begin
        if (!resetN) begin
            RGBout <= 8'h00;
        end else begin
            RGBout <= TRANSPARENT_ENCODING;

            if (InsideRectangle) begin
                RGBout <= object_colors[offsetY][offsetX];
            end
        end
    end

    assign drawingRequest = (RGBout != TRANSPARENT_ENCODING);

endmodule