module	claw_bitmap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 6;  // 2^6 = 64 
localparam  int OBJECT_NUMBER_OF_X_BITS = 6;  // 2^6 = 64 


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

// claw bitmap

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h7C ;// RGB value in the bitmap representing a transparent pixel 

logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [7:0] object_colors = {
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h00,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h00,8'h00,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFA,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h71,8'h71,8'h71,8'h71,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'hF9,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hF9,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF9,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'hFF,8'hFF,8'hFF,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C},
	{8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C,8'h7C}
};

 
 
// pipeline (ff) to get the pixel color from the array 	 

//////////--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN)
		RGBout <=	8'h7C;

	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default  

		if (InsideRectangle == 1'b1 )
			RGBout <= object_colors[offsetY][offsetX]; 
	end
		
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING); // get optional transparent command from the bitmpap   

endmodule