 module circle_object      	
	(
   // Input, Output Ports
	input  logic [6:0] alpha, //degree between 0-90
	input  logic [2:0] shift_radius, // if the user wants a smaller pixel
	output logic [9:0] dx,
	output logic [9:0] dy
   );

localparam logic sine_loc = 1'b0;
localparam logic cosine_loc = 1'b1;

// the range is between 0-2048, first col is sine, second cosine
logic [9:0] degree_covnerter [0:90][0:1] = '{
'{10'd0, 10'd1023},
'{10'd18, 10'd1023},
'{10'd36, 10'd1023},
'{10'd54, 10'd1023},
'{10'd71, 10'd1022},
'{10'd89, 10'd1020},
'{10'd107, 10'd1018},
'{10'd125, 10'd1016},
'{10'd143, 10'd1014},
'{10'd160, 10'd1011},
'{10'd178, 10'd1008},
'{10'd195, 10'd1005},
'{10'd213, 10'd1002},
'{10'd230, 10'd998},
'{10'd248, 10'd994},
'{10'd265, 10'd989},
'{10'd282, 10'd984},
'{10'd299, 10'd979},
'{10'd316, 10'd974},
'{10'd333, 10'd968},
'{10'd350, 10'd962},
'{10'd367, 10'd956},
'{10'd384, 10'd949},
'{10'd400, 10'd943},
'{10'd416, 10'd935},
'{10'd433, 10'd928},
'{10'd449, 10'd920},
'{10'd465, 10'd912},
'{10'd481, 10'd904},
'{10'd496, 10'd896},
'{10'd512, 10'd887},
'{10'd527, 10'd878},
'{10'd543, 10'd868},
'{10'd558, 10'd859},
'{10'd573, 10'd849},
'{10'd587, 10'd839},
'{10'd602, 10'd828},
'{10'd616, 10'd818},
'{10'd630, 10'd807},
'{10'd644, 10'd796},
'{10'd658, 10'd784},
'{10'd672, 10'd773},
'{10'd685, 10'd761},
'{10'd698, 10'd749},
'{10'd711, 10'd737},
'{10'd724, 10'd724},
'{10'd737, 10'd711},
'{10'd749, 10'd698},
'{10'd761, 10'd685},
'{10'd773, 10'd672},
'{10'd784, 10'd658},
'{10'd796, 10'd644},
'{10'd807, 10'd630},
'{10'd818, 10'd616},
'{10'd828, 10'd602},
'{10'd839, 10'd587},
'{10'd849, 10'd573},
'{10'd859, 10'd558},
'{10'd868, 10'd543},
'{10'd878, 10'd527},
'{10'd887, 10'd512},
'{10'd896, 10'd496},
'{10'd904, 10'd481},
'{10'd912, 10'd465},
'{10'd920, 10'd449},
'{10'd928, 10'd433},
'{10'd935, 10'd416},
'{10'd943, 10'd400},
'{10'd949, 10'd384},
'{10'd956, 10'd367},
'{10'd962, 10'd350},
'{10'd968, 10'd333},
'{10'd974, 10'd316},
'{10'd979, 10'd299},
'{10'd984, 10'd282},
'{10'd989, 10'd265},
'{10'd994, 10'd248},
'{10'd998, 10'd230},
'{10'd1002, 10'd213},
'{10'd1005, 10'd195},
'{10'd1008, 10'd178},
'{10'd1011, 10'd160},
'{10'd1014, 10'd143},
'{10'd1016, 10'd125},
'{10'd1018, 10'd107},
'{10'd1020, 10'd89},
'{10'd1022, 10'd71},
'{10'd1023, 10'd54},
'{10'd1023, 10'd36},
'{10'd1023, 10'd18},
'{10'd1023, 10'd0}
};


always_comb begin
	dx = degree_covnerter[alpha][cosine_loc] >> shift_radius;
	dy = degree_covnerter[alpha][sine_loc] >> shift_radius;
	if (alpha > 7'd90) begin
		dx = degree_covnerter[7'd90][cosine_loc] >> shift_radius;
		dy = degree_covnerter[7'd90][sine_loc] >> shift_radius;
	end
end
	
endmodule